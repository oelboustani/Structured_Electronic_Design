"CS Stage - Drive"
* C:\Users\maboa\Desktop\Structured Electronic Design\slicap\examples\Active Antenna\CS_stage_Drive\cir\CSstage_Drive.asc
M1 N001 V_GS 0 0 C18nmos l={L} w={W} m={m}
E1 V_GS 0 N003 0 1k
V1 N001 N003 {V_DS}
I1 0 N003 {I_DS}
M2 N002 In 0 0 C18nmos l={L} w={W} ad={w*500n} as={w*500n} pd={2*w+1u} ps={2*w+1u} m={m}
E2 In N004 V_GS 0 1
V2 N002 Out {V_DS}
I2 0 Out {I_DS}
R1 Out 0 {R_L}
V3 N005 0 AC 1
C2 N005 N004 {C_s}
.param L=180n W=40u M=6 I_DS=7m V_DS=0.4
.op
.lib CMOS18TT.lib
;op
.param R_L=50 C_s=1.5p
.ac dec 10 1k 100G
.backanno
.end
