"Drive"
* C:\Users\Tom\OneDrive\Desktop\Assignments\Q2\Structured Eelectronic Design\Assignment3_reorganised\Assignment 3\Drive.asc
M3 N004 N002 N001 N001 C18pmos l=180n w=40u m=11
M4 N004 N006 N005 N005 C18nmos l=180n w=40u m=3
V1 N001 0 0.9
V2 0 N005 0.9
R2 out N004 50
R3 0 out 50
V4 N003 N006 {V_d_bias/2}
V3 N003 0 SINE(0 300m 30meg)
C1 N004 0 2.5p
V5 N002 N003 {V_d_bias/2}
.param V_B=0.3 V_d_bias=0.66
.lib CMOS18TT.lib
;dc V3 -0.5 0.5 0.01
.step param V_B 0 0.5 0.05
.meas DC Ibias FIND (I(V1)+I(V2))/2 AT 0
.tran 0 50n 0 100p
.backanno
.end
